module selectPC(
    input wire ;

    output wire [63:0] predPC_o;
);



endmodule