module updatePC (
    input wire icode_i;
    input wire cnd;
    input wire [63:0] valC;

    output wire[63:0] PC
);
    
endmodule